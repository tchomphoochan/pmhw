////////////////////////////////////////////////////////////////////////////////
//  Filename      : Puppet.bsv
//  Description   : Execution unit for Puppetmaster.
////////////////////////////////////////////////////////////////////////////////
import PmCore::*;
import PmIfc::*;

////////////////////////////////////////////////////////////////////////////////
/// Module interface.
////////////////////////////////////////////////////////////////////////////////
typedef 5 LogTransactionDelayBase;

typedef TExp#(LogTransactionDelayBase) TransactionDelayBase;

typedef Bit#(TAdd#(LogTransactionObjectCount, LogTransactionDelayBase)) TransactionTimer;

interface Puppet;
    method Action start(RenamedTransaction tr);
    method Bool isDone();
endinterface

////////////////////////////////////////////////////////////////////////////////
/// Numeric constants.
////////////////////////////////////////////////////////////////////////////////
Integer delayBase = valueOf(TransactionDelayBase);

////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////
///
/// Puppet implementation.
///
/// Simulates executing a transaction by waiting for a number of cycles. This
/// number is calculated by multiplying TransactionDelayBase by the number of
/// objects (total, not distinct) in the transaction.
///
////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////
module mkPuppet(Puppet);
    ////////////////////////////////////////////////////////////////////////////////
    /// Design elements.
    ////////////////////////////////////////////////////////////////////////////////
    Reg#(TransactionTimer) timeLeft[2] <- mkCReg(2, 0);

    ////////////////////////////////////////////////////////////////////////////////
    /// Rules.
    ////////////////////////////////////////////////////////////////////////////////
    (* no_implicit_conditions, fire_when_enabled *)
    rule incTime if (0 < timeLeft[0]);
        timeLeft[0] <= timeLeft[0] - 1;
    endrule

    ////////////////////////////////////////////////////////////////////////////////
    /// Interface connections and methods.
    ////////////////////////////////////////////////////////////////////////////////
    method Action start(RenamedTransaction tr);
        let objCount = tr.readObjectCount + tr.writtenObjectCount;
        timeLeft[1] <= extend(objCount) * fromInteger(delayBase);
    endmethod

    method Bool isDone();
        return timeLeft[1] == 0;
    endmethod
endmodule
