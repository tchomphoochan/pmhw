typedef 1024 NumberLiveObjects;
typedef Bit#(NumberLiveObjects) ObjectSet;

typedef 16 SizeSchedulingPool;
typedef Bit#(SizeSchedulingPool) TransactionIds;
