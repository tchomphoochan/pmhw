typedef 10 LogNumberLiveObjects;
typedef 3 LogSizeRenamerBuffer;
typedef 3 LogNumberShards;
typedef 3 LogNumberHashes;
typedef 3 LogSizeSchedulingPool;
typedef 1 LogNumberComparators;
typedef 3 LogNumberPuppets;
