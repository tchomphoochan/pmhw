typedef 2 LogNumberRenamerThreads;
typedef 2 LogNumberShards;
typedef 6 LogSizeShard;
typedef 6 LogNumberHashes;
typedef 1 LogNumberComparators;
typedef 1 LogNumberSchedulingRounds;
typedef 3 LogNumberPuppets;
typedef 6 NumberAddressOffsetBits;
typedef 7 LogSizeRenamerBuffer;

/* Values for golden tests
typedef 3 LogNumberRenamerThreads;
typedef 3 LogNumberShards;
typedef 7 LogSizeShard;
typedef 4 LogNumberHashes;
typedef 1 LogNumberComparators;
typedef 1 LogNumberSchedulingRounds;
typedef 3 LogNumberPuppets;
typedef 6 NumberAddressOffsetBits;
typedef 3 LogSizeRenamerBuffer;
*/