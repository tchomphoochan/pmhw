typedef 10 LogNumberLiveObjects;
typedef TExp#(LogNumberLiveObjects) NumberLiveObjects;
typedef Bit#(NumberLiveObjects) ObjectSet;

typedef 4 LogSizeSchedulingPool;
typedef TExp#(LogSizeSchedulingPool) SizeSchedulingPool;
typedef Bit#(SizeSchedulingPool) TransactionIds;