typedef 3 LogNumberRenamerThreads;
typedef 3 LogNumberShards;
typedef 7 LogSizeShard;
typedef 4 LogNumberHashes;
typedef 1 LogNumberComparators;
typedef 1 LogNumberSchedulingRounds;
typedef 3 LogNumberPuppets;
typedef 6 NumberAddressOffsetBits;
typedef 8 LogSizeRenamerBuffer;
