////////////////////////////////////////////////////////////////////////////////
//  Filename      : Puppet.bsv
//  Description   : Execution unit for Puppetmaster.
////////////////////////////////////////////////////////////////////////////////
import PmCore::*;
import PmIfc::*;

////////////////////////////////////////////////////////////////////////////////
/// Module interface.
////////////////////////////////////////////////////////////////////////////////
interface Puppet;
    method Action start(RenamedTransaction tr);
    method Bool isDone();
endinterface

////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////
///
/// Puppet implementation.
///
/// Simulates executing a transaction by waiting for a number of cycles. This
/// number is calculated by multiplying TransactionDelayBase by the number of
/// objects (total, not distinct) in the transaction.
///
////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////
(* synthesize *)
module mkPuppet(Puppet);
    ////////////////////////////////////////////////////////////////////////////////
    /// Design elements.
    ////////////////////////////////////////////////////////////////////////////////
    Reg#(Timestamp) timeLeft[2] <- mkCReg(2, 0);

    ////////////////////////////////////////////////////////////////////////////////
    /// Rules.
    ////////////////////////////////////////////////////////////////////////////////
    (* no_implicit_conditions, fire_when_enabled *)
    rule incTime if (0 < timeLeft[0]);
        timeLeft[0] <= timeLeft[0] - 1;
    endrule

    ////////////////////////////////////////////////////////////////////////////////
    /// Interface connections and methods.
    ////////////////////////////////////////////////////////////////////////////////
    method Action start(RenamedTransaction tr);
        Timestamp trDuration = case (tr.trType) matches
            DatabaseRead : 2000;
            DatabaseWrite : 2000;
            DatabaseIncrement : 4000;
            DatabaseSwap : 8000;
            MessageFetch : 1800;
            MessagePost : 240;
        endcase;
        timeLeft[1] <= trDuration;
    endmethod

    method Bool isDone();
        return timeLeft[1] == 0;
    endmethod
endmodule
